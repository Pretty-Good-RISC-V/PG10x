interface DebugModule;
endinterface

module mkDebugModule(DebugModule);
endmodule
