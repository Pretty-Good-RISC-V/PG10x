typedef 1 FetchStageNumber;
typedef 2 DecodeStageNumber;
typedef 3 ExecutionStageNumber;
typedef 4 MemoryAccessStageNumber;
typedef 5 WritebackStageNumber;